module simple_wire();



endmodule
