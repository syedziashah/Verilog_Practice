module tb_simple_wire();



endmodule
